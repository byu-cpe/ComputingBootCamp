module top(
  input LIOB33_X0Y11_IOB_X0Y11_IPAD,
  input RIOB33_X43Y25_IOB_X1Y26_IPAD,
  output LIOB33_X0Y19_IOB_X0Y19_OPAD,
  output LIOB33_X0Y19_IOB_X0Y20_OPAD,
  output LIOB33_X0Y3_IOB_X0Y3_OPAD,
  output LIOB33_X0Y43_IOB_X0Y43_OPAD
  );
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A5Q;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_AMUX;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_AO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_AO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_AQ;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_A_XOR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B5Q;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_BMUX;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_BO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_BO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_BQ;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_B_XOR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_CLK;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_CO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_CO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_C_XOR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_DO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_DO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_D_XOR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X0Y19_SR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_AO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_AO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_A_XOR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_BO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_BO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_B_XOR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_CO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_CO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_C_XOR;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D1;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D2;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D3;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D4;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_DO5;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_DO6;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D_CY;
  wire [0:0] CLBLL_L_X2Y19_SLICE_X1Y19_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_A5_FDRE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(1'b1),
.D(CLBLL_L_X2Y19_SLICE_X0Y19_AO5),
.Q(CLBLL_L_X2Y19_SLICE_X0Y19_A5Q),
.R(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_B5_FDRE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(1'b1),
.D(CLBLL_L_X2Y19_SLICE_X0Y19_BO5),
.Q(CLBLL_L_X2Y19_SLICE_X0Y19_B5Q),
.R(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_A_FDRE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(1'b1),
.D(CLBLL_L_X2Y19_SLICE_X0Y19_AO6),
.Q(CLBLL_L_X2Y19_SLICE_X0Y19_AQ),
.R(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_B_FDRE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(1'b1),
.D(CLBLL_L_X2Y19_SLICE_X0Y19_BO6),
.Q(CLBLL_L_X2Y19_SLICE_X0Y19_BQ),
.R(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'b0000111100001111000011110000111100111100001111000011110000111100)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y19_SLICE_X0Y19_A5Q),
.I2(CLBLL_L_X2Y19_SLICE_X0Y19_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X0Y19_AO5),
.O6(CLBLL_L_X2Y19_SLICE_X0Y19_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'b0011110000111100110011001100110001101010011010101010101010101010)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_BLUT (
.I0(CLBLL_L_X2Y19_SLICE_X0Y19_B5Q),
.I1(CLBLL_L_X2Y19_SLICE_X0Y19_BQ),
.I2(CLBLL_L_X2Y19_SLICE_X0Y19_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y19_SLICE_X0Y19_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X0Y19_BO5),
.O6(CLBLL_L_X2Y19_SLICE_X0Y19_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'b0000000000000000000000000000000000000000000000000000000000000000)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X0Y19_CO5),
.O6(CLBLL_L_X2Y19_SLICE_X0Y19_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'b0000000000000000000000000000000000000000000000000000000000000000)
  ) CLBLL_L_X2Y19_SLICE_X0Y19_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X0Y19_DO5),
.O6(CLBLL_L_X2Y19_SLICE_X0Y19_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'b0000000000000000000000000000000000000000000000000000000000000000)
  ) CLBLL_L_X2Y19_SLICE_X1Y19_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X1Y19_AO5),
.O6(CLBLL_L_X2Y19_SLICE_X1Y19_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'b0000000000000000000000000000000000000000000000000000000000000000)
  ) CLBLL_L_X2Y19_SLICE_X1Y19_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X1Y19_BO5),
.O6(CLBLL_L_X2Y19_SLICE_X1Y19_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'b0000000000000000000000000000000000000000000000000000000000000000)
  ) CLBLL_L_X2Y19_SLICE_X1Y19_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X1Y19_CO5),
.O6(CLBLL_L_X2Y19_SLICE_X1Y19_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'b0000000000000000000000000000000000000000000000000000000000000000)
  ) CLBLL_L_X2Y19_SLICE_X1Y19_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y19_SLICE_X1Y19_DO5),
.O6(CLBLL_L_X2Y19_SLICE_X1Y19_DO6)
  );


  (* KEEP, DONT_TOUCH *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O)
  );


  (* KEEP, DONT_TOUCH *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUF (
.I(CLBLL_L_X2Y19_SLICE_X0Y19_AQ),
.O(LIOB33_X0Y3_IOB_X0Y3_OPAD)
  );


  (* KEEP, DONT_TOUCH *)
  IBUF #(
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(LIOB33_X0Y11_IOB_X0Y11_IPAD),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y19_OBUF (
.I(CLBLL_L_X2Y19_SLICE_X0Y19_B5Q),
.O(LIOB33_X0Y19_IOB_X0Y19_OPAD)
  );


  (* KEEP, DONT_TOUCH *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y20_OBUF (
.I(CLBLL_L_X2Y19_SLICE_X0Y19_BQ),
.O(LIOB33_X0Y19_IOB_X0Y20_OPAD)
  );


  (* KEEP, DONT_TOUCH *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(CLBLL_L_X2Y19_SLICE_X0Y19_A5Q),
.O(LIOB33_X0Y43_IOB_X0Y43_OPAD)
  );


  (* KEEP, DONT_TOUCH *)
  IBUF #(
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(RIOB33_X43Y25_IOB_X1Y26_IPAD),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );
  assign CLBLL_L_X2Y19_SLICE_X0Y19_A = CLBLL_L_X2Y19_SLICE_X0Y19_AO6;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_B = CLBLL_L_X2Y19_SLICE_X0Y19_BO6;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_C = CLBLL_L_X2Y19_SLICE_X0Y19_CO6;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_D = CLBLL_L_X2Y19_SLICE_X0Y19_DO6;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_AMUX = CLBLL_L_X2Y19_SLICE_X0Y19_A5Q;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_BMUX = CLBLL_L_X2Y19_SLICE_X0Y19_B5Q;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_A = CLBLL_L_X2Y19_SLICE_X1Y19_AO6;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_B = CLBLL_L_X2Y19_SLICE_X1Y19_BO6;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_C = CLBLL_L_X2Y19_SLICE_X1Y19_CO6;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_D = CLBLL_L_X2Y19_SLICE_X1Y19_DO6;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOI3_X0Y11_ILOGIC_X0Y11_D;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ = LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ = LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ = LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ = LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ = LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOI3_X43Y25_ILOGIC_X1Y26_D;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_D3 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_D4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_D5 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  assign LIOB33_X0Y19_IOB_X0Y20_O = CLBLL_L_X2Y19_SLICE_X0Y19_BQ;
  assign LIOB33_X0Y19_IOB_X0Y19_O = CLBLL_L_X2Y19_SLICE_X0Y19_B5Q;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_A1 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_A2 = CLBLL_L_X2Y19_SLICE_X0Y19_A5Q;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_A3 = CLBLL_L_X2Y19_SLICE_X0Y19_AQ;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_A4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_A5 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_A6 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_B1 = CLBLL_L_X2Y19_SLICE_X0Y19_B5Q;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_B2 = CLBLL_L_X2Y19_SLICE_X0Y19_BQ;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_B3 = CLBLL_L_X2Y19_SLICE_X0Y19_AQ;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_B4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_B5 = CLBLL_L_X2Y19_SLICE_X0Y19_A5Q;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_B6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_C1 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_C2 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_C3 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_C4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_C5 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_C6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y3_O = CLBLL_L_X2Y19_SLICE_X0Y19_AQ;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_D1 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_D2 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_D3 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_D4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_D5 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_D6 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X0Y19_SR = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOB33_X0Y43_IOB_X0Y43_O = CLBLL_L_X2Y19_SLICE_X0Y19_A5Q;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_A1 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_A2 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_A3 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_A4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_A5 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_A6 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_B1 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_B2 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_B3 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_B4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_B5 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_B6 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_C1 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_C2 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_C3 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_C4 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_C5 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_C6 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_D1 = 1'b1;
  assign CLBLL_L_X2Y19_SLICE_X1Y19_D2 = 1'b1;
endmodule